** Profile: "SCHEMATIC1-Components Sweep"  [ C:\Users\kpapa01\Desktop\NYU POLY\SEMESTERS\NYU SPRING 13\EE3114 Fundamentals of Electronics I\OrCad Capture CIS Demo\HW 00\EE3114 Hwk0 Resistor Divider-PSpiceFiles\SCHEMATIC1\Components Sweep.sim ] 

** Creating circuit file "Components Sweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\OrCAD\OrCAD_16.3_Demo\tools\PSpice\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.DC LIN PARAM Rval 1k 10k 1k 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
