** Profile: "SCHEMATIC1-HW04 MOSFET"  [ C:\Users\kpapa01\Desktop\NYU POLY\SEMESTERS\NYU SPRING 13\EE3114 Fundamentals of Electronics I\HW\HW04 MOSFET-PSpiceFiles\SCHEMATIC1\HW04 MOSFET.sim ] 

** Creating circuit file "HW04 MOSFET.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\OrCAD\OrCAD_16.3_Demo\tools\PSpice\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 25msec 0 0.001msec 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
